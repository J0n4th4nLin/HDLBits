module top_module(output zero);
    
    //// Module body starts after semicolon
    assign zero = 1'b0;

endmodule
/*
    This question requires the output to be 0.
        So the right side of b is 0.
*/